// ECE423_QSYS.v

// Generated using ACDS version 15.1 193

`timescale 1 ps / 1 ps
module ECE423_QSYS (
	);

	ECE423_QSYS_QSYS_0 qsys_0 (
	);

endmodule
