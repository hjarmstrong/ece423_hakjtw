// ECE423_QSYS_QSYS_0.v

// Generated using ACDS version 15.1 193

`timescale 1 ps / 1 ps
module ECE423_QSYS_QSYS_0 (
	);

	ECE423_QSYS_QSYS_0_QSYS_0 qsys_0 (
	);

endmodule
